module re_e200(input clk);
endmodule
