module re_e200();
endmodule
